// TODO
// instantiate letter select here
module morse_code_detector(..);

